---------------------------------------------------------------------------
-- (c) Copyright: OscillatorIMP Digital
-- Author : Gwenhael Goavec-Merou<gwenhael.goavec-merou@trabucayre.com>
-- Creation date : 2015/04/08
---------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.ALL;

entity nco_counter_cos_rom_a12_d16 is
port (
	clk : in std_logic;
	addr_a : in std_logic_vector(11 downto 0);
	addr_b : in std_logic_vector(11 downto 0);
	data_a : out std_logic_vector(15 downto 0);
	data_b : out std_logic_vector(15 downto 0));
end entity nco_counter_cos_rom_a12_d16;

architecture behavioral of nco_counter_cos_rom_a12_d16 is

	signal i: integer range 0 to 2**12-1 :=0;
	type mem is array ( 0 to 2**12-1) of 
			std_logic_vector(15 downto 0);

	constant my_Rom : mem := (
		"0111111111111111",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111101",
		"0111111111111101",
		"0111111111111100",
		"0111111111111011",
		"0111111111111011",
		"0111111111111010",
		"0111111111111001",
		"0111111111111000",
		"0111111111110111",
		"0111111111110110",
		"0111111111110101",
		"0111111111110011",
		"0111111111110010",
		"0111111111110001",
		"0111111111101111",
		"0111111111101110",
		"0111111111101100",
		"0111111111101010",
		"0111111111101000",
		"0111111111100110",
		"0111111111100100",
		"0111111111100010",
		"0111111111100000",
		"0111111111011110",
		"0111111111011100",
		"0111111111011001",
		"0111111111010111",
		"0111111111010101",
		"0111111111010010",
		"0111111111001111",
		"0111111111001101",
		"0111111111001010",
		"0111111111000111",
		"0111111111000100",
		"0111111111000001",
		"0111111110111110",
		"0111111110111011",
		"0111111110110111",
		"0111111110110100",
		"0111111110110000",
		"0111111110101101",
		"0111111110101001",
		"0111111110100110",
		"0111111110100010",
		"0111111110011110",
		"0111111110011010",
		"0111111110010110",
		"0111111110010010",
		"0111111110001110",
		"0111111110001010",
		"0111111110000110",
		"0111111110000001",
		"0111111101111101",
		"0111111101111000",
		"0111111101110100",
		"0111111101101111",
		"0111111101101010",
		"0111111101100110",
		"0111111101100001",
		"0111111101011100",
		"0111111101010111",
		"0111111101010010",
		"0111111101001100",
		"0111111101000111",
		"0111111101000010",
		"0111111100111100",
		"0111111100110111",
		"0111111100110001",
		"0111111100101100",
		"0111111100100110",
		"0111111100100000",
		"0111111100011010",
		"0111111100010100",
		"0111111100001110",
		"0111111100001000",
		"0111111100000010",
		"0111111011111100",
		"0111111011110101",
		"0111111011101111",
		"0111111011101000",
		"0111111011100010",
		"0111111011011011",
		"0111111011010100",
		"0111111011001110",
		"0111111011000111",
		"0111111011000000",
		"0111111010111001",
		"0111111010110010",
		"0111111010101010",
		"0111111010100011",
		"0111111010011100",
		"0111111010010100",
		"0111111010001101",
		"0111111010000101",
		"0111111001111110",
		"0111111001110110",
		"0111111001101110",
		"0111111001100110",
		"0111111001011110",
		"0111111001010110",
		"0111111001001110",
		"0111111001000110",
		"0111111000111110",
		"0111111000110110",
		"0111111000101101",
		"0111111000100101",
		"0111111000011100",
		"0111111000010011",
		"0111111000001011",
		"0111111000000010",
		"0111110111111001",
		"0111110111110000",
		"0111110111100111",
		"0111110111011110",
		"0111110111010101",
		"0111110111001100",
		"0111110111000010",
		"0111110110111001",
		"0111110110110000",
		"0111110110100110",
		"0111110110011100",
		"0111110110010011",
		"0111110110001001",
		"0111110101111111",
		"0111110101110101",
		"0111110101101011",
		"0111110101100001",
		"0111110101010111",
		"0111110101001101",
		"0111110101000010",
		"0111110100111000",
		"0111110100101110",
		"0111110100100011",
		"0111110100011000",
		"0111110100001110",
		"0111110100000011",
		"0111110011111000",
		"0111110011101101",
		"0111110011100010",
		"0111110011010111",
		"0111110011001100",
		"0111110011000001",
		"0111110010110110",
		"0111110010101010",
		"0111110010011111",
		"0111110010010011",
		"0111110010001000",
		"0111110001111100",
		"0111110001110000",
		"0111110001100101",
		"0111110001011001",
		"0111110001001101",
		"0111110001000001",
		"0111110000110101",
		"0111110000101001",
		"0111110000011100",
		"0111110000010000",
		"0111110000000100",
		"0111101111110111",
		"0111101111101011",
		"0111101111011110",
		"0111101111010001",
		"0111101111000100",
		"0111101110111000",
		"0111101110101011",
		"0111101110011110",
		"0111101110010001",
		"0111101110000011",
		"0111101101110110",
		"0111101101101001",
		"0111101101011100",
		"0111101101001110",
		"0111101101000001",
		"0111101100110011",
		"0111101100100101",
		"0111101100011000",
		"0111101100001010",
		"0111101011111100",
		"0111101011101110",
		"0111101011100000",
		"0111101011010010",
		"0111101011000100",
		"0111101010110101",
		"0111101010100111",
		"0111101010011001",
		"0111101010001010",
		"0111101001111100",
		"0111101001101101",
		"0111101001011110",
		"0111101001001111",
		"0111101001000001",
		"0111101000110010",
		"0111101000100011",
		"0111101000010100",
		"0111101000000100",
		"0111100111110101",
		"0111100111100110",
		"0111100111010111",
		"0111100111000111",
		"0111100110111000",
		"0111100110101000",
		"0111100110011000",
		"0111100110001001",
		"0111100101111001",
		"0111100101101001",
		"0111100101011001",
		"0111100101001001",
		"0111100100111001",
		"0111100100101001",
		"0111100100011001",
		"0111100100001000",
		"0111100011111000",
		"0111100011100111",
		"0111100011010111",
		"0111100011000110",
		"0111100010110110",
		"0111100010100101",
		"0111100010010100",
		"0111100010000011",
		"0111100001110010",
		"0111100001100001",
		"0111100001010000",
		"0111100000111111",
		"0111100000101110",
		"0111100000011100",
		"0111100000001011",
		"0111011111111001",
		"0111011111101000",
		"0111011111010110",
		"0111011111000100",
		"0111011110110011",
		"0111011110100001",
		"0111011110001111",
		"0111011101111101",
		"0111011101101011",
		"0111011101011001",
		"0111011101000111",
		"0111011100110100",
		"0111011100100010",
		"0111011100010000",
		"0111011011111101",
		"0111011011101010",
		"0111011011011000",
		"0111011011000101",
		"0111011010110010",
		"0111011010100000",
		"0111011010001101",
		"0111011001111010",
		"0111011001100111",
		"0111011001010011",
		"0111011001000000",
		"0111011000101101",
		"0111011000011010",
		"0111011000000110",
		"0111010111110011",
		"0111010111011111",
		"0111010111001100",
		"0111010110111000",
		"0111010110100100",
		"0111010110010000",
		"0111010101111100",
		"0111010101101000",
		"0111010101010100",
		"0111010101000000",
		"0111010100101100",
		"0111010100011000",
		"0111010100000011",
		"0111010011101111",
		"0111010011011011",
		"0111010011000110",
		"0111010010110001",
		"0111010010011101",
		"0111010010001000",
		"0111010001110011",
		"0111010001011110",
		"0111010001001001",
		"0111010000110100",
		"0111010000011111",
		"0111010000001010",
		"0111001111110101",
		"0111001111011111",
		"0111001111001010",
		"0111001110110101",
		"0111001110011111",
		"0111001110001001",
		"0111001101110100",
		"0111001101011110",
		"0111001101001000",
		"0111001100110010",
		"0111001100011100",
		"0111001100000110",
		"0111001011110000",
		"0111001011011010",
		"0111001011000100",
		"0111001010101110",
		"0111001010010111",
		"0111001010000001",
		"0111001001101010",
		"0111001001010100",
		"0111001000111101",
		"0111001000100110",
		"0111001000010000",
		"0111000111111001",
		"0111000111100010",
		"0111000111001011",
		"0111000110110100",
		"0111000110011101",
		"0111000110000110",
		"0111000101101110",
		"0111000101010111",
		"0111000101000000",
		"0111000100101000",
		"0111000100010001",
		"0111000011111001",
		"0111000011100001",
		"0111000011001010",
		"0111000010110010",
		"0111000010011010",
		"0111000010000010",
		"0111000001101010",
		"0111000001010010",
		"0111000000111010",
		"0111000000100010",
		"0111000000001001",
		"0110111111110001",
		"0110111111011001",
		"0110111111000000",
		"0110111110101000",
		"0110111110001111",
		"0110111101110110",
		"0110111101011110",
		"0110111101000101",
		"0110111100101100",
		"0110111100010011",
		"0110111011111010",
		"0110111011100001",
		"0110111011001000",
		"0110111010101111",
		"0110111010010101",
		"0110111001111100",
		"0110111001100011",
		"0110111001001001",
		"0110111000110000",
		"0110111000010110",
		"0110110111111100",
		"0110110111100011",
		"0110110111001001",
		"0110110110101111",
		"0110110110010101",
		"0110110101111011",
		"0110110101100001",
		"0110110101000111",
		"0110110100101100",
		"0110110100010010",
		"0110110011111000",
		"0110110011011101",
		"0110110011000011",
		"0110110010101000",
		"0110110010001110",
		"0110110001110011",
		"0110110001011000",
		"0110110000111110",
		"0110110000100011",
		"0110110000001000",
		"0110101111101101",
		"0110101111010010",
		"0110101110110111",
		"0110101110011100",
		"0110101110000000",
		"0110101101100101",
		"0110101101001010",
		"0110101100101110",
		"0110101100010011",
		"0110101011110111",
		"0110101011011011",
		"0110101011000000",
		"0110101010100100",
		"0110101010001000",
		"0110101001101100",
		"0110101001010000",
		"0110101000110100",
		"0110101000011000",
		"0110100111111100",
		"0110100111100000",
		"0110100111000100",
		"0110100110100111",
		"0110100110001011",
		"0110100101101110",
		"0110100101010010",
		"0110100100110101",
		"0110100100011001",
		"0110100011111100",
		"0110100011011111",
		"0110100011000010",
		"0110100010100101",
		"0110100010001000",
		"0110100001101011",
		"0110100001001110",
		"0110100000110001",
		"0110100000010100",
		"0110011111110111",
		"0110011111011001",
		"0110011110111100",
		"0110011110011110",
		"0110011110000001",
		"0110011101100011",
		"0110011101000101",
		"0110011100101000",
		"0110011100001010",
		"0110011011101100",
		"0110011011001110",
		"0110011010110000",
		"0110011010010010",
		"0110011001110100",
		"0110011001010110",
		"0110011000111000",
		"0110011000011001",
		"0110010111111011",
		"0110010111011101",
		"0110010110111110",
		"0110010110100000",
		"0110010110000001",
		"0110010101100010",
		"0110010101000100",
		"0110010100100101",
		"0110010100000110",
		"0110010011100111",
		"0110010011001000",
		"0110010010101001",
		"0110010010001010",
		"0110010001101011",
		"0110010001001100",
		"0110010000101101",
		"0110010000001101",
		"0110001111101110",
		"0110001111001110",
		"0110001110101111",
		"0110001110001111",
		"0110001101110000",
		"0110001101010000",
		"0110001100110000",
		"0110001100010001",
		"0110001011110001",
		"0110001011010001",
		"0110001010110001",
		"0110001010010001",
		"0110001001110001",
		"0110001001010001",
		"0110001000110000",
		"0110001000010000",
		"0110000111110000",
		"0110000111001111",
		"0110000110101111",
		"0110000110001110",
		"0110000101101110",
		"0110000101001101",
		"0110000100101101",
		"0110000100001100",
		"0110000011101011",
		"0110000011001010",
		"0110000010101001",
		"0110000010001000",
		"0110000001100111",
		"0110000001000110",
		"0110000000100101",
		"0110000000000100",
		"0101111111100010",
		"0101111111000001",
		"0101111110100000",
		"0101111101111110",
		"0101111101011101",
		"0101111100111011",
		"0101111100011010",
		"0101111011111000",
		"0101111011010110",
		"0101111010110100",
		"0101111010010011",
		"0101111001110001",
		"0101111001001111",
		"0101111000101101",
		"0101111000001011",
		"0101110111101001",
		"0101110111000110",
		"0101110110100100",
		"0101110110000010",
		"0101110101011111",
		"0101110100111101",
		"0101110100011011",
		"0101110011111000",
		"0101110011010110",
		"0101110010110011",
		"0101110010010000",
		"0101110001101101",
		"0101110001001011",
		"0101110000101000",
		"0101110000000101",
		"0101101111100010",
		"0101101110111111",
		"0101101110011100",
		"0101101101111001",
		"0101101101010110",
		"0101101100110010",
		"0101101100001111",
		"0101101011101100",
		"0101101011001000",
		"0101101010100101",
		"0101101010000001",
		"0101101001011110",
		"0101101000111010",
		"0101101000010110",
		"0101100111110011",
		"0101100111001111",
		"0101100110101011",
		"0101100110000111",
		"0101100101100011",
		"0101100100111111",
		"0101100100011011",
		"0101100011110111",
		"0101100011010011",
		"0101100010101111",
		"0101100010001010",
		"0101100001100110",
		"0101100001000010",
		"0101100000011101",
		"0101011111111001",
		"0101011111010100",
		"0101011110110000",
		"0101011110001011",
		"0101011101100110",
		"0101011101000010",
		"0101011100011101",
		"0101011011111000",
		"0101011011010011",
		"0101011010101110",
		"0101011010001001",
		"0101011001100100",
		"0101011000111111",
		"0101011000011010",
		"0101010111110100",
		"0101010111001111",
		"0101010110101010",
		"0101010110000101",
		"0101010101011111",
		"0101010100111010",
		"0101010100010100",
		"0101010011101111",
		"0101010011001001",
		"0101010010100011",
		"0101010001111101",
		"0101010001011000",
		"0101010000110010",
		"0101010000001100",
		"0101001111100110",
		"0101001111000000",
		"0101001110011010",
		"0101001101110100",
		"0101001101001110",
		"0101001100101000",
		"0101001100000001",
		"0101001011011011",
		"0101001010110101",
		"0101001010001110",
		"0101001001101000",
		"0101001001000001",
		"0101001000011011",
		"0101000111110100",
		"0101000111001110",
		"0101000110100111",
		"0101000110000000",
		"0101000101011001",
		"0101000100110011",
		"0101000100001100",
		"0101000011100101",
		"0101000010111110",
		"0101000010010111",
		"0101000001110000",
		"0101000001001001",
		"0101000000100001",
		"0100111111111010",
		"0100111111010011",
		"0100111110101100",
		"0100111110000100",
		"0100111101011101",
		"0100111100110101",
		"0100111100001110",
		"0100111011100110",
		"0100111010111111",
		"0100111010010111",
		"0100111001101111",
		"0100111001001000",
		"0100111000100000",
		"0100110111111000",
		"0100110111010000",
		"0100110110101000",
		"0100110110000000",
		"0100110101011000",
		"0100110100110000",
		"0100110100001000",
		"0100110011100000",
		"0100110010111000",
		"0100110010001111",
		"0100110001100111",
		"0100110000111111",
		"0100110000010110",
		"0100101111101110",
		"0100101111000101",
		"0100101110011101",
		"0100101101110100",
		"0100101101001100",
		"0100101100100011",
		"0100101011111010",
		"0100101011010010",
		"0100101010101001",
		"0100101010000000",
		"0100101001010111",
		"0100101000101110",
		"0100101000000101",
		"0100100111011100",
		"0100100110110011",
		"0100100110001010",
		"0100100101100001",
		"0100100100111000",
		"0100100100001110",
		"0100100011100101",
		"0100100010111100",
		"0100100010010010",
		"0100100001101001",
		"0100100000111111",
		"0100100000010110",
		"0100011111101100",
		"0100011111000011",
		"0100011110011001",
		"0100011101101111",
		"0100011101000110",
		"0100011100011100",
		"0100011011110010",
		"0100011011001000",
		"0100011010011110",
		"0100011001110100",
		"0100011001001010",
		"0100011000100000",
		"0100010111110110",
		"0100010111001100",
		"0100010110100010",
		"0100010101111000",
		"0100010101001110",
		"0100010100100011",
		"0100010011111001",
		"0100010011001111",
		"0100010010100100",
		"0100010001111010",
		"0100010001001111",
		"0100010000100101",
		"0100001111111010",
		"0100001111010000",
		"0100001110100101",
		"0100001101111010",
		"0100001101010000",
		"0100001100100101",
		"0100001011111010",
		"0100001011001111",
		"0100001010100100",
		"0100001001111001",
		"0100001001001110",
		"0100001000100011",
		"0100000111111000",
		"0100000111001101",
		"0100000110100010",
		"0100000101110111",
		"0100000101001100",
		"0100000100100000",
		"0100000011110101",
		"0100000011001010",
		"0100000010011110",
		"0100000001110011",
		"0100000001000111",
		"0100000000011100",
		"0011111111110000",
		"0011111111000101",
		"0011111110011001",
		"0011111101101110",
		"0011111101000010",
		"0011111100010110",
		"0011111011101011",
		"0011111010111111",
		"0011111010010011",
		"0011111001100111",
		"0011111000111011",
		"0011111000001111",
		"0011110111100011",
		"0011110110110111",
		"0011110110001011",
		"0011110101011111",
		"0011110100110011",
		"0011110100000111",
		"0011110011011011",
		"0011110010101110",
		"0011110010000010",
		"0011110001010110",
		"0011110000101001",
		"0011101111111101",
		"0011101111010001",
		"0011101110100100",
		"0011101101111000",
		"0011101101001011",
		"0011101100011111",
		"0011101011110010",
		"0011101011000101",
		"0011101010011001",
		"0011101001101100",
		"0011101000111111",
		"0011101000010010",
		"0011100111100110",
		"0011100110111001",
		"0011100110001100",
		"0011100101011111",
		"0011100100110010",
		"0011100100000101",
		"0011100011011000",
		"0011100010101011",
		"0011100001111110",
		"0011100001010001",
		"0011100000100100",
		"0011011111110110",
		"0011011111001001",
		"0011011110011100",
		"0011011101101111",
		"0011011101000001",
		"0011011100010100",
		"0011011011100111",
		"0011011010111001",
		"0011011010001100",
		"0011011001011110",
		"0011011000110001",
		"0011011000000011",
		"0011010111010110",
		"0011010110101000",
		"0011010101111010",
		"0011010101001101",
		"0011010100011111",
		"0011010011110001",
		"0011010011000011",
		"0011010010010110",
		"0011010001101000",
		"0011010000111010",
		"0011010000001100",
		"0011001111011110",
		"0011001110110000",
		"0011001110000010",
		"0011001101010100",
		"0011001100100110",
		"0011001011111000",
		"0011001011001010",
		"0011001010011100",
		"0011001001101101",
		"0011001000111111",
		"0011001000010001",
		"0011000111100011",
		"0011000110110100",
		"0011000110000110",
		"0011000101011000",
		"0011000100101001",
		"0011000011111011",
		"0011000011001100",
		"0011000010011110",
		"0011000001101111",
		"0011000001000001",
		"0011000000010010",
		"0010111111100100",
		"0010111110110101",
		"0010111110000110",
		"0010111101011000",
		"0010111100101001",
		"0010111011111010",
		"0010111011001100",
		"0010111010011101",
		"0010111001101110",
		"0010111000111111",
		"0010111000010000",
		"0010110111100001",
		"0010110110110010",
		"0010110110000011",
		"0010110101010100",
		"0010110100100101",
		"0010110011110110",
		"0010110011000111",
		"0010110010011000",
		"0010110001101001",
		"0010110000111010",
		"0010110000001011",
		"0010101111011011",
		"0010101110101100",
		"0010101101111101",
		"0010101101001110",
		"0010101100011110",
		"0010101011101111",
		"0010101011000000",
		"0010101010010000",
		"0010101001100001",
		"0010101000110001",
		"0010101000000010",
		"0010100111010010",
		"0010100110100011",
		"0010100101110011",
		"0010100101000100",
		"0010100100010100",
		"0010100011100101",
		"0010100010110101",
		"0010100010000101",
		"0010100001010110",
		"0010100000100110",
		"0010011111110110",
		"0010011111000110",
		"0010011110010111",
		"0010011101100111",
		"0010011100110111",
		"0010011100000111",
		"0010011011010111",
		"0010011010100111",
		"0010011001110111",
		"0010011001000111",
		"0010011000010111",
		"0010010111100111",
		"0010010110110111",
		"0010010110000111",
		"0010010101010111",
		"0010010100100111",
		"0010010011110111",
		"0010010011000111",
		"0010010010010111",
		"0010010001100111",
		"0010010000110110",
		"0010010000000110",
		"0010001111010110",
		"0010001110100110",
		"0010001101110101",
		"0010001101000101",
		"0010001100010101",
		"0010001011100100",
		"0010001010110100",
		"0010001010000100",
		"0010001001010011",
		"0010001000100011",
		"0010000111110010",
		"0010000111000010",
		"0010000110010001",
		"0010000101100001",
		"0010000100110000",
		"0010000100000000",
		"0010000011001111",
		"0010000010011111",
		"0010000001101110",
		"0010000000111101",
		"0010000000001101",
		"0001111111011100",
		"0001111110101011",
		"0001111101111011",
		"0001111101001010",
		"0001111100011001",
		"0001111011101000",
		"0001111010111000",
		"0001111010000111",
		"0001111001010110",
		"0001111000100101",
		"0001110111110100",
		"0001110111000011",
		"0001110110010011",
		"0001110101100010",
		"0001110100110001",
		"0001110100000000",
		"0001110011001111",
		"0001110010011110",
		"0001110001101101",
		"0001110000111100",
		"0001110000001011",
		"0001101111011010",
		"0001101110101001",
		"0001101101111000",
		"0001101101000110",
		"0001101100010101",
		"0001101011100100",
		"0001101010110011",
		"0001101010000010",
		"0001101001010001",
		"0001101000100000",
		"0001100111101110",
		"0001100110111101",
		"0001100110001100",
		"0001100101011011",
		"0001100100101001",
		"0001100011111000",
		"0001100011000111",
		"0001100010010101",
		"0001100001100100",
		"0001100000110011",
		"0001100000000001",
		"0001011111010000",
		"0001011110011111",
		"0001011101101101",
		"0001011100111100",
		"0001011100001010",
		"0001011011011001",
		"0001011010100111",
		"0001011001110110",
		"0001011001000100",
		"0001011000010011",
		"0001010111100001",
		"0001010110110000",
		"0001010101111110",
		"0001010101001101",
		"0001010100011011",
		"0001010011101010",
		"0001010010111000",
		"0001010010000110",
		"0001010001010101",
		"0001010000100011",
		"0001001111110010",
		"0001001111000000",
		"0001001110001110",
		"0001001101011101",
		"0001001100101011",
		"0001001011111001",
		"0001001011000111",
		"0001001010010110",
		"0001001001100100",
		"0001001000110010",
		"0001001000000000",
		"0001000111001111",
		"0001000110011101",
		"0001000101101011",
		"0001000100111001",
		"0001000100000111",
		"0001000011010110",
		"0001000010100100",
		"0001000001110010",
		"0001000001000000",
		"0001000000001110",
		"0000111111011100",
		"0000111110101011",
		"0000111101111001",
		"0000111101000111",
		"0000111100010101",
		"0000111011100011",
		"0000111010110001",
		"0000111001111111",
		"0000111001001101",
		"0000111000011011",
		"0000110111101001",
		"0000110110110111",
		"0000110110000101",
		"0000110101010011",
		"0000110100100001",
		"0000110011101111",
		"0000110010111101",
		"0000110010001011",
		"0000110001011001",
		"0000110000100111",
		"0000101111110101",
		"0000101111000011",
		"0000101110010001",
		"0000101101011111",
		"0000101100101101",
		"0000101011111011",
		"0000101011001001",
		"0000101010010111",
		"0000101001100101",
		"0000101000110010",
		"0000101000000000",
		"0000100111001110",
		"0000100110011100",
		"0000100101101010",
		"0000100100111000",
		"0000100100000110",
		"0000100011010100",
		"0000100010100001",
		"0000100001101111",
		"0000100000111101",
		"0000100000001011",
		"0000011111011001",
		"0000011110100111",
		"0000011101110100",
		"0000011101000010",
		"0000011100010000",
		"0000011011011110",
		"0000011010101100",
		"0000011001111010",
		"0000011001000111",
		"0000011000010101",
		"0000010111100011",
		"0000010110110001",
		"0000010101111110",
		"0000010101001100",
		"0000010100011010",
		"0000010011101000",
		"0000010010110110",
		"0000010010000011",
		"0000010001010001",
		"0000010000011111",
		"0000001111101101",
		"0000001110111010",
		"0000001110001000",
		"0000001101010110",
		"0000001100100100",
		"0000001011110001",
		"0000001010111111",
		"0000001010001101",
		"0000001001011011",
		"0000001000101000",
		"0000000111110110",
		"0000000111000100",
		"0000000110010010",
		"0000000101011111",
		"0000000100101101",
		"0000000011111011",
		"0000000011001001",
		"0000000010010110",
		"0000000001100100",
		"0000000000110010",
		"0000000000000000",
		"1111111111001110",
		"1111111110011100",
		"1111111101101010",
		"1111111100110111",
		"1111111100000101",
		"1111111011010011",
		"1111111010100001",
		"1111111001101110",
		"1111111000111100",
		"1111111000001010",
		"1111110111011000",
		"1111110110100101",
		"1111110101110011",
		"1111110101000001",
		"1111110100001111",
		"1111110011011100",
		"1111110010101010",
		"1111110001111000",
		"1111110001000110",
		"1111110000010011",
		"1111101111100001",
		"1111101110101111",
		"1111101101111101",
		"1111101101001010",
		"1111101100011000",
		"1111101011100110",
		"1111101010110100",
		"1111101010000010",
		"1111101001001111",
		"1111101000011101",
		"1111100111101011",
		"1111100110111001",
		"1111100110000110",
		"1111100101010100",
		"1111100100100010",
		"1111100011110000",
		"1111100010111110",
		"1111100010001100",
		"1111100001011001",
		"1111100000100111",
		"1111011111110101",
		"1111011111000011",
		"1111011110010001",
		"1111011101011111",
		"1111011100101100",
		"1111011011111010",
		"1111011011001000",
		"1111011010010110",
		"1111011001100100",
		"1111011000110010",
		"1111011000000000",
		"1111010111001110",
		"1111010110011011",
		"1111010101101001",
		"1111010100110111",
		"1111010100000101",
		"1111010011010011",
		"1111010010100001",
		"1111010001101111",
		"1111010000111101",
		"1111010000001011",
		"1111001111011001",
		"1111001110100111",
		"1111001101110101",
		"1111001101000011",
		"1111001100010001",
		"1111001011011111",
		"1111001010101101",
		"1111001001111011",
		"1111001001001001",
		"1111001000010111",
		"1111000111100101",
		"1111000110110011",
		"1111000110000001",
		"1111000101001111",
		"1111000100011101",
		"1111000011101011",
		"1111000010111001",
		"1111000010000111",
		"1111000001010101",
		"1111000000100100",
		"1110111111110010",
		"1110111111000000",
		"1110111110001110",
		"1110111101011100",
		"1110111100101010",
		"1110111011111001",
		"1110111011000111",
		"1110111010010101",
		"1110111001100011",
		"1110111000110001",
		"1110111000000000",
		"1110110111001110",
		"1110110110011100",
		"1110110101101010",
		"1110110100111001",
		"1110110100000111",
		"1110110011010101",
		"1110110010100011",
		"1110110001110010",
		"1110110001000000",
		"1110110000001110",
		"1110101111011101",
		"1110101110101011",
		"1110101101111010",
		"1110101101001000",
		"1110101100010110",
		"1110101011100101",
		"1110101010110011",
		"1110101010000010",
		"1110101001010000",
		"1110101000011111",
		"1110100111101101",
		"1110100110111100",
		"1110100110001010",
		"1110100101011001",
		"1110100100100111",
		"1110100011110110",
		"1110100011000100",
		"1110100010010011",
		"1110100001100001",
		"1110100000110000",
		"1110011111111111",
		"1110011111001101",
		"1110011110011100",
		"1110011101101011",
		"1110011100111001",
		"1110011100001000",
		"1110011011010111",
		"1110011010100101",
		"1110011001110100",
		"1110011001000011",
		"1110011000010010",
		"1110010111100000",
		"1110010110101111",
		"1110010101111110",
		"1110010101001101",
		"1110010100011100",
		"1110010011101011",
		"1110010010111010",
		"1110010010001000",
		"1110010001010111",
		"1110010000100110",
		"1110001111110101",
		"1110001111000100",
		"1110001110010011",
		"1110001101100010",
		"1110001100110001",
		"1110001100000000",
		"1110001011001111",
		"1110001010011110",
		"1110001001101101",
		"1110001000111101",
		"1110001000001100",
		"1110000111011011",
		"1110000110101010",
		"1110000101111001",
		"1110000101001000",
		"1110000100011000",
		"1110000011100111",
		"1110000010110110",
		"1110000010000101",
		"1110000001010101",
		"1110000000100100",
		"1101111111110011",
		"1101111111000011",
		"1101111110010010",
		"1101111101100001",
		"1101111100110001",
		"1101111100000000",
		"1101111011010000",
		"1101111010011111",
		"1101111001101111",
		"1101111000111110",
		"1101111000001110",
		"1101110111011101",
		"1101110110101101",
		"1101110101111100",
		"1101110101001100",
		"1101110100011100",
		"1101110011101011",
		"1101110010111011",
		"1101110010001011",
		"1101110001011010",
		"1101110000101010",
		"1101101111111010",
		"1101101111001010",
		"1101101110011001",
		"1101101101101001",
		"1101101100111001",
		"1101101100001001",
		"1101101011011001",
		"1101101010101001",
		"1101101001111001",
		"1101101001001001",
		"1101101000011001",
		"1101100111101001",
		"1101100110111001",
		"1101100110001001",
		"1101100101011001",
		"1101100100101001",
		"1101100011111001",
		"1101100011001001",
		"1101100010011001",
		"1101100001101001",
		"1101100000111010",
		"1101100000001010",
		"1101011111011010",
		"1101011110101010",
		"1101011101111011",
		"1101011101001011",
		"1101011100011011",
		"1101011011101100",
		"1101011010111100",
		"1101011010001101",
		"1101011001011101",
		"1101011000101110",
		"1101010111111110",
		"1101010111001111",
		"1101010110011111",
		"1101010101110000",
		"1101010101000000",
		"1101010100010001",
		"1101010011100010",
		"1101010010110010",
		"1101010010000011",
		"1101010001010100",
		"1101010000100101",
		"1101001111110101",
		"1101001111000110",
		"1101001110010111",
		"1101001101101000",
		"1101001100111001",
		"1101001100001010",
		"1101001011011011",
		"1101001010101100",
		"1101001001111101",
		"1101001001001110",
		"1101001000011111",
		"1101000111110000",
		"1101000111000001",
		"1101000110010010",
		"1101000101100011",
		"1101000100110100",
		"1101000100000110",
		"1101000011010111",
		"1101000010101000",
		"1101000001111010",
		"1101000001001011",
		"1101000000011100",
		"1100111111101110",
		"1100111110111111",
		"1100111110010001",
		"1100111101100010",
		"1100111100110100",
		"1100111100000101",
		"1100111011010111",
		"1100111010101000",
		"1100111001111010",
		"1100111001001100",
		"1100111000011101",
		"1100110111101111",
		"1100110111000001",
		"1100110110010011",
		"1100110101100100",
		"1100110100110110",
		"1100110100001000",
		"1100110011011010",
		"1100110010101100",
		"1100110001111110",
		"1100110001010000",
		"1100110000100010",
		"1100101111110100",
		"1100101111000110",
		"1100101110011000",
		"1100101101101010",
		"1100101100111101",
		"1100101100001111",
		"1100101011100001",
		"1100101010110011",
		"1100101010000110",
		"1100101001011000",
		"1100101000101010",
		"1100100111111101",
		"1100100111001111",
		"1100100110100010",
		"1100100101110100",
		"1100100101000111",
		"1100100100011001",
		"1100100011101100",
		"1100100010111111",
		"1100100010010001",
		"1100100001100100",
		"1100100000110111",
		"1100100000001010",
		"1100011111011100",
		"1100011110101111",
		"1100011110000010",
		"1100011101010101",
		"1100011100101000",
		"1100011011111011",
		"1100011011001110",
		"1100011010100001",
		"1100011001110100",
		"1100011001000111",
		"1100011000011010",
		"1100010111101110",
		"1100010111000001",
		"1100010110010100",
		"1100010101100111",
		"1100010100111011",
		"1100010100001110",
		"1100010011100001",
		"1100010010110101",
		"1100010010001000",
		"1100010001011100",
		"1100010000101111",
		"1100010000000011",
		"1100001111010111",
		"1100001110101010",
		"1100001101111110",
		"1100001101010010",
		"1100001100100101",
		"1100001011111001",
		"1100001011001101",
		"1100001010100001",
		"1100001001110101",
		"1100001001001001",
		"1100001000011101",
		"1100000111110001",
		"1100000111000101",
		"1100000110011001",
		"1100000101101101",
		"1100000101000001",
		"1100000100010101",
		"1100000011101010",
		"1100000010111110",
		"1100000010010010",
		"1100000001100111",
		"1100000000111011",
		"1100000000010000",
		"1011111111100100",
		"1011111110111001",
		"1011111110001101",
		"1011111101100010",
		"1011111100110110",
		"1011111100001011",
		"1011111011100000",
		"1011111010110100",
		"1011111010001001",
		"1011111001011110",
		"1011111000110011",
		"1011111000001000",
		"1011110111011101",
		"1011110110110010",
		"1011110110000111",
		"1011110101011100",
		"1011110100110001",
		"1011110100000110",
		"1011110011011011",
		"1011110010110000",
		"1011110010000110",
		"1011110001011011",
		"1011110000110000",
		"1011110000000110",
		"1011101111011011",
		"1011101110110001",
		"1011101110000110",
		"1011101101011100",
		"1011101100110001",
		"1011101100000111",
		"1011101011011101",
		"1011101010110010",
		"1011101010001000",
		"1011101001011110",
		"1011101000110100",
		"1011101000001010",
		"1011100111100000",
		"1011100110110110",
		"1011100110001100",
		"1011100101100010",
		"1011100100111000",
		"1011100100001110",
		"1011100011100100",
		"1011100010111010",
		"1011100010010001",
		"1011100001100111",
		"1011100000111101",
		"1011100000010100",
		"1011011111101010",
		"1011011111000001",
		"1011011110010111",
		"1011011101101110",
		"1011011101000100",
		"1011011100011011",
		"1011011011110010",
		"1011011011001000",
		"1011011010011111",
		"1011011001110110",
		"1011011001001101",
		"1011011000100100",
		"1011010111111011",
		"1011010111010010",
		"1011010110101001",
		"1011010110000000",
		"1011010101010111",
		"1011010100101110",
		"1011010100000110",
		"1011010011011101",
		"1011010010110100",
		"1011010010001100",
		"1011010001100011",
		"1011010000111011",
		"1011010000010010",
		"1011001111101010",
		"1011001111000001",
		"1011001110011001",
		"1011001101110001",
		"1011001101001000",
		"1011001100100000",
		"1011001011111000",
		"1011001011010000",
		"1011001010101000",
		"1011001010000000",
		"1011001001011000",
		"1011001000110000",
		"1011001000001000",
		"1011000111100000",
		"1011000110111000",
		"1011000110010001",
		"1011000101101001",
		"1011000101000001",
		"1011000100011010",
		"1011000011110010",
		"1011000011001011",
		"1011000010100011",
		"1011000001111100",
		"1011000001010100",
		"1011000000101101",
		"1011000000000110",
		"1010111111011111",
		"1010111110110111",
		"1010111110010000",
		"1010111101101001",
		"1010111101000010",
		"1010111100011011",
		"1010111011110100",
		"1010111011001101",
		"1010111010100111",
		"1010111010000000",
		"1010111001011001",
		"1010111000110010",
		"1010111000001100",
		"1010110111100101",
		"1010110110111111",
		"1010110110011000",
		"1010110101110010",
		"1010110101001011",
		"1010110100100101",
		"1010110011111111",
		"1010110011011000",
		"1010110010110010",
		"1010110010001100",
		"1010110001100110",
		"1010110001000000",
		"1010110000011010",
		"1010101111110100",
		"1010101111001110",
		"1010101110101000",
		"1010101110000011",
		"1010101101011101",
		"1010101100110111",
		"1010101100010001",
		"1010101011101100",
		"1010101011000110",
		"1010101010100001",
		"1010101001111011",
		"1010101001010110",
		"1010101000110001",
		"1010101000001100",
		"1010100111100110",
		"1010100111000001",
		"1010100110011100",
		"1010100101110111",
		"1010100101010010",
		"1010100100101101",
		"1010100100001000",
		"1010100011100011",
		"1010100010111110",
		"1010100010011010",
		"1010100001110101",
		"1010100001010000",
		"1010100000101100",
		"1010100000000111",
		"1010011111100011",
		"1010011110111110",
		"1010011110011010",
		"1010011101110110",
		"1010011101010001",
		"1010011100101101",
		"1010011100001001",
		"1010011011100101",
		"1010011011000001",
		"1010011010011101",
		"1010011001111001",
		"1010011001010101",
		"1010011000110001",
		"1010011000001101",
		"1010010111101010",
		"1010010111000110",
		"1010010110100010",
		"1010010101111111",
		"1010010101011011",
		"1010010100111000",
		"1010010100010100",
		"1010010011110001",
		"1010010011001110",
		"1010010010101010",
		"1010010010000111",
		"1010010001100100",
		"1010010001000001",
		"1010010000011110",
		"1010001111111011",
		"1010001111011000",
		"1010001110110101",
		"1010001110010011",
		"1010001101110000",
		"1010001101001101",
		"1010001100101010",
		"1010001100001000",
		"1010001011100101",
		"1010001011000011",
		"1010001010100001",
		"1010001001111110",
		"1010001001011100",
		"1010001000111010",
		"1010001000010111",
		"1010000111110101",
		"1010000111010011",
		"1010000110110001",
		"1010000110001111",
		"1010000101101101",
		"1010000101001100",
		"1010000100101010",
		"1010000100001000",
		"1010000011100110",
		"1010000011000101",
		"1010000010100011",
		"1010000010000010",
		"1010000001100000",
		"1010000000111111",
		"1010000000011110",
		"1001111111111100",
		"1001111111011011",
		"1001111110111010",
		"1001111110011001",
		"1001111101111000",
		"1001111101010111",
		"1001111100110110",
		"1001111100010101",
		"1001111011110100",
		"1001111011010011",
		"1001111010110011",
		"1001111010010010",
		"1001111001110010",
		"1001111001010001",
		"1001111000110001",
		"1001111000010000",
		"1001110111110000",
		"1001110111010000",
		"1001110110101111",
		"1001110110001111",
		"1001110101101111",
		"1001110101001111",
		"1001110100101111",
		"1001110100001111",
		"1001110011101111",
		"1001110011010000",
		"1001110010110000",
		"1001110010010000",
		"1001110001110001",
		"1001110001010001",
		"1001110000110010",
		"1001110000010010",
		"1001101111110011",
		"1001101111010011",
		"1001101110110100",
		"1001101110010101",
		"1001101101110110",
		"1001101101010111",
		"1001101100111000",
		"1001101100011001",
		"1001101011111010",
		"1001101011011011",
		"1001101010111100",
		"1001101010011110",
		"1001101001111111",
		"1001101001100000",
		"1001101001000010",
		"1001101000100011",
		"1001101000000101",
		"1001100111100111",
		"1001100111001000",
		"1001100110101010",
		"1001100110001100",
		"1001100101101110",
		"1001100101010000",
		"1001100100110010",
		"1001100100010100",
		"1001100011110110",
		"1001100011011000",
		"1001100010111011",
		"1001100010011101",
		"1001100001111111",
		"1001100001100010",
		"1001100001000100",
		"1001100000100111",
		"1001100000001001",
		"1001011111101100",
		"1001011111001111",
		"1001011110110010",
		"1001011110010101",
		"1001011101111000",
		"1001011101011011",
		"1001011100111110",
		"1001011100100001",
		"1001011100000100",
		"1001011011100111",
		"1001011011001011",
		"1001011010101110",
		"1001011010010010",
		"1001011001110101",
		"1001011001011001",
		"1001011000111100",
		"1001011000100000",
		"1001011000000100",
		"1001010111101000",
		"1001010111001100",
		"1001010110110000",
		"1001010110010100",
		"1001010101111000",
		"1001010101011100",
		"1001010101000000",
		"1001010100100101",
		"1001010100001001",
		"1001010011101101",
		"1001010011010010",
		"1001010010110110",
		"1001010010011011",
		"1001010010000000",
		"1001010001100100",
		"1001010001001001",
		"1001010000101110",
		"1001010000010011",
		"1001001111111000",
		"1001001111011101",
		"1001001111000010",
		"1001001110101000",
		"1001001110001101",
		"1001001101110010",
		"1001001101011000",
		"1001001100111101",
		"1001001100100011",
		"1001001100001000",
		"1001001011101110",
		"1001001011010100",
		"1001001010111001",
		"1001001010011111",
		"1001001010000101",
		"1001001001101011",
		"1001001001010001",
		"1001001000110111",
		"1001001000011101",
		"1001001000000100",
		"1001000111101010",
		"1001000111010000",
		"1001000110110111",
		"1001000110011101",
		"1001000110000100",
		"1001000101101011",
		"1001000101010001",
		"1001000100111000",
		"1001000100011111",
		"1001000100000110",
		"1001000011101101",
		"1001000011010100",
		"1001000010111011",
		"1001000010100010",
		"1001000010001010",
		"1001000001110001",
		"1001000001011000",
		"1001000001000000",
		"1001000000100111",
		"1001000000001111",
		"1000111111110111",
		"1000111111011110",
		"1000111111000110",
		"1000111110101110",
		"1000111110010110",
		"1000111101111110",
		"1000111101100110",
		"1000111101001110",
		"1000111100110110",
		"1000111100011111",
		"1000111100000111",
		"1000111011101111",
		"1000111011011000",
		"1000111011000000",
		"1000111010101001",
		"1000111010010010",
		"1000111001111010",
		"1000111001100011",
		"1000111001001100",
		"1000111000110101",
		"1000111000011110",
		"1000111000000111",
		"1000110111110000",
		"1000110111011010",
		"1000110111000011",
		"1000110110101100",
		"1000110110010110",
		"1000110101111111",
		"1000110101101001",
		"1000110101010010",
		"1000110100111100",
		"1000110100100110",
		"1000110100010000",
		"1000110011111010",
		"1000110011100100",
		"1000110011001110",
		"1000110010111000",
		"1000110010100010",
		"1000110010001100",
		"1000110001110111",
		"1000110001100001",
		"1000110001001011",
		"1000110000110110",
		"1000110000100001",
		"1000110000001011",
		"1000101111110110",
		"1000101111100001",
		"1000101111001100",
		"1000101110110111",
		"1000101110100010",
		"1000101110001101",
		"1000101101111000",
		"1000101101100011",
		"1000101101001111",
		"1000101100111010",
		"1000101100100101",
		"1000101100010001",
		"1000101011111101",
		"1000101011101000",
		"1000101011010100",
		"1000101011000000",
		"1000101010101100",
		"1000101010011000",
		"1000101010000100",
		"1000101001110000",
		"1000101001011100",
		"1000101001001000",
		"1000101000110100",
		"1000101000100001",
		"1000101000001101",
		"1000100111111010",
		"1000100111100110",
		"1000100111010011",
		"1000100111000000",
		"1000100110101101",
		"1000100110011001",
		"1000100110000110",
		"1000100101110011",
		"1000100101100000",
		"1000100101001110",
		"1000100100111011",
		"1000100100101000",
		"1000100100010110",
		"1000100100000011",
		"1000100011110000",
		"1000100011011110",
		"1000100011001100",
		"1000100010111001",
		"1000100010100111",
		"1000100010010101",
		"1000100010000011",
		"1000100001110001",
		"1000100001011111",
		"1000100001001101",
		"1000100000111100",
		"1000100000101010",
		"1000100000011000",
		"1000100000000111",
		"1000011111110101",
		"1000011111100100",
		"1000011111010010",
		"1000011111000001",
		"1000011110110000",
		"1000011110011111",
		"1000011110001110",
		"1000011101111101",
		"1000011101101100",
		"1000011101011011",
		"1000011101001010",
		"1000011100111010",
		"1000011100101001",
		"1000011100011001",
		"1000011100001000",
		"1000011011111000",
		"1000011011100111",
		"1000011011010111",
		"1000011011000111",
		"1000011010110111",
		"1000011010100111",
		"1000011010010111",
		"1000011010000111",
		"1000011001110111",
		"1000011001101000",
		"1000011001011000",
		"1000011001001000",
		"1000011000111001",
		"1000011000101001",
		"1000011000011010",
		"1000011000001011",
		"1000010111111100",
		"1000010111101100",
		"1000010111011101",
		"1000010111001110",
		"1000010110111111",
		"1000010110110001",
		"1000010110100010",
		"1000010110010011",
		"1000010110000100",
		"1000010101110110",
		"1000010101100111",
		"1000010101011001",
		"1000010101001011",
		"1000010100111100",
		"1000010100101110",
		"1000010100100000",
		"1000010100010010",
		"1000010100000100",
		"1000010011110110",
		"1000010011101000",
		"1000010011011011",
		"1000010011001101",
		"1000010010111111",
		"1000010010110010",
		"1000010010100100",
		"1000010010010111",
		"1000010010001010",
		"1000010001111101",
		"1000010001101111",
		"1000010001100010",
		"1000010001010101",
		"1000010001001000",
		"1000010000111100",
		"1000010000101111",
		"1000010000100010",
		"1000010000010101",
		"1000010000001001",
		"1000001111111100",
		"1000001111110000",
		"1000001111100100",
		"1000001111010111",
		"1000001111001011",
		"1000001110111111",
		"1000001110110011",
		"1000001110100111",
		"1000001110011011",
		"1000001110010000",
		"1000001110000100",
		"1000001101111000",
		"1000001101101101",
		"1000001101100001",
		"1000001101010110",
		"1000001101001010",
		"1000001100111111",
		"1000001100110100",
		"1000001100101001",
		"1000001100011110",
		"1000001100010011",
		"1000001100001000",
		"1000001011111101",
		"1000001011110010",
		"1000001011101000",
		"1000001011011101",
		"1000001011010010",
		"1000001011001000",
		"1000001010111110",
		"1000001010110011",
		"1000001010101001",
		"1000001010011111",
		"1000001010010101",
		"1000001010001011",
		"1000001010000001",
		"1000001001110111",
		"1000001001101101",
		"1000001001100100",
		"1000001001011010",
		"1000001001010000",
		"1000001001000111",
		"1000001000111110",
		"1000001000110100",
		"1000001000101011",
		"1000001000100010",
		"1000001000011001",
		"1000001000010000",
		"1000001000000111",
		"1000000111111110",
		"1000000111110101",
		"1000000111101101",
		"1000000111100100",
		"1000000111011011",
		"1000000111010011",
		"1000000111001010",
		"1000000111000010",
		"1000000110111010",
		"1000000110110010",
		"1000000110101010",
		"1000000110100010",
		"1000000110011010",
		"1000000110010010",
		"1000000110001010",
		"1000000110000010",
		"1000000101111011",
		"1000000101110011",
		"1000000101101100",
		"1000000101100100",
		"1000000101011101",
		"1000000101010110",
		"1000000101001110",
		"1000000101000111",
		"1000000101000000",
		"1000000100111001",
		"1000000100110010",
		"1000000100101100",
		"1000000100100101",
		"1000000100011110",
		"1000000100011000",
		"1000000100010001",
		"1000000100001011",
		"1000000100000100",
		"1000000011111110",
		"1000000011111000",
		"1000000011110010",
		"1000000011101100",
		"1000000011100110",
		"1000000011100000",
		"1000000011011010",
		"1000000011010100",
		"1000000011001111",
		"1000000011001001",
		"1000000011000100",
		"1000000010111110",
		"1000000010111001",
		"1000000010110100",
		"1000000010101110",
		"1000000010101001",
		"1000000010100100",
		"1000000010011111",
		"1000000010011010",
		"1000000010010110",
		"1000000010010001",
		"1000000010001100",
		"1000000010001000",
		"1000000010000011",
		"1000000001111111",
		"1000000001111010",
		"1000000001110110",
		"1000000001110010",
		"1000000001101110",
		"1000000001101010",
		"1000000001100110",
		"1000000001100010",
		"1000000001011110",
		"1000000001011010",
		"1000000001010111",
		"1000000001010011",
		"1000000001010000",
		"1000000001001100",
		"1000000001001001",
		"1000000001000101",
		"1000000001000010",
		"1000000000111111",
		"1000000000111100",
		"1000000000111001",
		"1000000000110110",
		"1000000000110011",
		"1000000000110001",
		"1000000000101110",
		"1000000000101011",
		"1000000000101001",
		"1000000000100111",
		"1000000000100100",
		"1000000000100010",
		"1000000000100000",
		"1000000000011110",
		"1000000000011100",
		"1000000000011010",
		"1000000000011000",
		"1000000000010110",
		"1000000000010100",
		"1000000000010010",
		"1000000000010001",
		"1000000000001111",
		"1000000000001110",
		"1000000000001101",
		"1000000000001011",
		"1000000000001010",
		"1000000000001001",
		"1000000000001000",
		"1000000000000111",
		"1000000000000110",
		"1000000000000101",
		"1000000000000101",
		"1000000000000100",
		"1000000000000011",
		"1000000000000011",
		"1000000000000010",
		"1000000000000010",
		"1000000000000010",
		"1000000000000010",
		"1000000000000010",
		"1000000000000001",
		"1000000000000010",
		"1000000000000010",
		"1000000000000010",
		"1000000000000010",
		"1000000000000010",
		"1000000000000011",
		"1000000000000011",
		"1000000000000100",
		"1000000000000101",
		"1000000000000101",
		"1000000000000110",
		"1000000000000111",
		"1000000000001000",
		"1000000000001001",
		"1000000000001010",
		"1000000000001011",
		"1000000000001101",
		"1000000000001110",
		"1000000000001111",
		"1000000000010001",
		"1000000000010010",
		"1000000000010100",
		"1000000000010110",
		"1000000000011000",
		"1000000000011010",
		"1000000000011100",
		"1000000000011110",
		"1000000000100000",
		"1000000000100010",
		"1000000000100100",
		"1000000000100111",
		"1000000000101001",
		"1000000000101011",
		"1000000000101110",
		"1000000000110001",
		"1000000000110011",
		"1000000000110110",
		"1000000000111001",
		"1000000000111100",
		"1000000000111111",
		"1000000001000010",
		"1000000001000101",
		"1000000001001001",
		"1000000001001100",
		"1000000001010000",
		"1000000001010011",
		"1000000001010111",
		"1000000001011010",
		"1000000001011110",
		"1000000001100010",
		"1000000001100110",
		"1000000001101010",
		"1000000001101110",
		"1000000001110010",
		"1000000001110110",
		"1000000001111010",
		"1000000001111111",
		"1000000010000011",
		"1000000010001000",
		"1000000010001100",
		"1000000010010001",
		"1000000010010110",
		"1000000010011010",
		"1000000010011111",
		"1000000010100100",
		"1000000010101001",
		"1000000010101110",
		"1000000010110100",
		"1000000010111001",
		"1000000010111110",
		"1000000011000100",
		"1000000011001001",
		"1000000011001111",
		"1000000011010100",
		"1000000011011010",
		"1000000011100000",
		"1000000011100110",
		"1000000011101100",
		"1000000011110010",
		"1000000011111000",
		"1000000011111110",
		"1000000100000100",
		"1000000100001011",
		"1000000100010001",
		"1000000100011000",
		"1000000100011110",
		"1000000100100101",
		"1000000100101100",
		"1000000100110010",
		"1000000100111001",
		"1000000101000000",
		"1000000101000111",
		"1000000101001110",
		"1000000101010110",
		"1000000101011101",
		"1000000101100100",
		"1000000101101100",
		"1000000101110011",
		"1000000101111011",
		"1000000110000010",
		"1000000110001010",
		"1000000110010010",
		"1000000110011010",
		"1000000110100010",
		"1000000110101010",
		"1000000110110010",
		"1000000110111010",
		"1000000111000010",
		"1000000111001010",
		"1000000111010011",
		"1000000111011011",
		"1000000111100100",
		"1000000111101101",
		"1000000111110101",
		"1000000111111110",
		"1000001000000111",
		"1000001000010000",
		"1000001000011001",
		"1000001000100010",
		"1000001000101011",
		"1000001000110100",
		"1000001000111110",
		"1000001001000111",
		"1000001001010000",
		"1000001001011010",
		"1000001001100100",
		"1000001001101101",
		"1000001001110111",
		"1000001010000001",
		"1000001010001011",
		"1000001010010101",
		"1000001010011111",
		"1000001010101001",
		"1000001010110011",
		"1000001010111110",
		"1000001011001000",
		"1000001011010010",
		"1000001011011101",
		"1000001011101000",
		"1000001011110010",
		"1000001011111101",
		"1000001100001000",
		"1000001100010011",
		"1000001100011110",
		"1000001100101001",
		"1000001100110100",
		"1000001100111111",
		"1000001101001010",
		"1000001101010110",
		"1000001101100001",
		"1000001101101101",
		"1000001101111000",
		"1000001110000100",
		"1000001110010000",
		"1000001110011011",
		"1000001110100111",
		"1000001110110011",
		"1000001110111111",
		"1000001111001011",
		"1000001111010111",
		"1000001111100100",
		"1000001111110000",
		"1000001111111100",
		"1000010000001001",
		"1000010000010101",
		"1000010000100010",
		"1000010000101111",
		"1000010000111100",
		"1000010001001000",
		"1000010001010101",
		"1000010001100010",
		"1000010001101111",
		"1000010001111101",
		"1000010010001010",
		"1000010010010111",
		"1000010010100100",
		"1000010010110010",
		"1000010010111111",
		"1000010011001101",
		"1000010011011011",
		"1000010011101000",
		"1000010011110110",
		"1000010100000100",
		"1000010100010010",
		"1000010100100000",
		"1000010100101110",
		"1000010100111100",
		"1000010101001011",
		"1000010101011001",
		"1000010101100111",
		"1000010101110110",
		"1000010110000100",
		"1000010110010011",
		"1000010110100010",
		"1000010110110001",
		"1000010110111111",
		"1000010111001110",
		"1000010111011101",
		"1000010111101100",
		"1000010111111100",
		"1000011000001011",
		"1000011000011010",
		"1000011000101001",
		"1000011000111001",
		"1000011001001000",
		"1000011001011000",
		"1000011001101000",
		"1000011001110111",
		"1000011010000111",
		"1000011010010111",
		"1000011010100111",
		"1000011010110111",
		"1000011011000111",
		"1000011011010111",
		"1000011011100111",
		"1000011011111000",
		"1000011100001000",
		"1000011100011001",
		"1000011100101001",
		"1000011100111010",
		"1000011101001010",
		"1000011101011011",
		"1000011101101100",
		"1000011101111101",
		"1000011110001110",
		"1000011110011111",
		"1000011110110000",
		"1000011111000001",
		"1000011111010010",
		"1000011111100100",
		"1000011111110101",
		"1000100000000111",
		"1000100000011000",
		"1000100000101010",
		"1000100000111100",
		"1000100001001101",
		"1000100001011111",
		"1000100001110001",
		"1000100010000011",
		"1000100010010101",
		"1000100010100111",
		"1000100010111001",
		"1000100011001100",
		"1000100011011110",
		"1000100011110000",
		"1000100100000011",
		"1000100100010110",
		"1000100100101000",
		"1000100100111011",
		"1000100101001110",
		"1000100101100000",
		"1000100101110011",
		"1000100110000110",
		"1000100110011001",
		"1000100110101101",
		"1000100111000000",
		"1000100111010011",
		"1000100111100110",
		"1000100111111010",
		"1000101000001101",
		"1000101000100001",
		"1000101000110100",
		"1000101001001000",
		"1000101001011100",
		"1000101001110000",
		"1000101010000100",
		"1000101010011000",
		"1000101010101100",
		"1000101011000000",
		"1000101011010100",
		"1000101011101000",
		"1000101011111101",
		"1000101100010001",
		"1000101100100101",
		"1000101100111010",
		"1000101101001111",
		"1000101101100011",
		"1000101101111000",
		"1000101110001101",
		"1000101110100010",
		"1000101110110111",
		"1000101111001100",
		"1000101111100001",
		"1000101111110110",
		"1000110000001011",
		"1000110000100001",
		"1000110000110110",
		"1000110001001011",
		"1000110001100001",
		"1000110001110111",
		"1000110010001100",
		"1000110010100010",
		"1000110010111000",
		"1000110011001110",
		"1000110011100100",
		"1000110011111010",
		"1000110100010000",
		"1000110100100110",
		"1000110100111100",
		"1000110101010010",
		"1000110101101001",
		"1000110101111111",
		"1000110110010110",
		"1000110110101100",
		"1000110111000011",
		"1000110111011010",
		"1000110111110000",
		"1000111000000111",
		"1000111000011110",
		"1000111000110101",
		"1000111001001100",
		"1000111001100011",
		"1000111001111010",
		"1000111010010010",
		"1000111010101001",
		"1000111011000000",
		"1000111011011000",
		"1000111011101111",
		"1000111100000111",
		"1000111100011111",
		"1000111100110110",
		"1000111101001110",
		"1000111101100110",
		"1000111101111110",
		"1000111110010110",
		"1000111110101110",
		"1000111111000110",
		"1000111111011110",
		"1000111111110111",
		"1001000000001111",
		"1001000000100111",
		"1001000001000000",
		"1001000001011000",
		"1001000001110001",
		"1001000010001010",
		"1001000010100010",
		"1001000010111011",
		"1001000011010100",
		"1001000011101101",
		"1001000100000110",
		"1001000100011111",
		"1001000100111000",
		"1001000101010001",
		"1001000101101011",
		"1001000110000100",
		"1001000110011101",
		"1001000110110111",
		"1001000111010000",
		"1001000111101010",
		"1001001000000100",
		"1001001000011101",
		"1001001000110111",
		"1001001001010001",
		"1001001001101011",
		"1001001010000101",
		"1001001010011111",
		"1001001010111001",
		"1001001011010100",
		"1001001011101110",
		"1001001100001000",
		"1001001100100011",
		"1001001100111101",
		"1001001101011000",
		"1001001101110010",
		"1001001110001101",
		"1001001110101000",
		"1001001111000010",
		"1001001111011101",
		"1001001111111000",
		"1001010000010011",
		"1001010000101110",
		"1001010001001001",
		"1001010001100100",
		"1001010010000000",
		"1001010010011011",
		"1001010010110110",
		"1001010011010010",
		"1001010011101101",
		"1001010100001001",
		"1001010100100101",
		"1001010101000000",
		"1001010101011100",
		"1001010101111000",
		"1001010110010100",
		"1001010110110000",
		"1001010111001100",
		"1001010111101000",
		"1001011000000100",
		"1001011000100000",
		"1001011000111100",
		"1001011001011001",
		"1001011001110101",
		"1001011010010010",
		"1001011010101110",
		"1001011011001011",
		"1001011011100111",
		"1001011100000100",
		"1001011100100001",
		"1001011100111110",
		"1001011101011011",
		"1001011101111000",
		"1001011110010101",
		"1001011110110010",
		"1001011111001111",
		"1001011111101100",
		"1001100000001001",
		"1001100000100111",
		"1001100001000100",
		"1001100001100010",
		"1001100001111111",
		"1001100010011101",
		"1001100010111011",
		"1001100011011000",
		"1001100011110110",
		"1001100100010100",
		"1001100100110010",
		"1001100101010000",
		"1001100101101110",
		"1001100110001100",
		"1001100110101010",
		"1001100111001000",
		"1001100111100111",
		"1001101000000101",
		"1001101000100011",
		"1001101001000010",
		"1001101001100000",
		"1001101001111111",
		"1001101010011110",
		"1001101010111100",
		"1001101011011011",
		"1001101011111010",
		"1001101100011001",
		"1001101100111000",
		"1001101101010111",
		"1001101101110110",
		"1001101110010101",
		"1001101110110100",
		"1001101111010011",
		"1001101111110011",
		"1001110000010010",
		"1001110000110010",
		"1001110001010001",
		"1001110001110001",
		"1001110010010000",
		"1001110010110000",
		"1001110011010000",
		"1001110011101111",
		"1001110100001111",
		"1001110100101111",
		"1001110101001111",
		"1001110101101111",
		"1001110110001111",
		"1001110110101111",
		"1001110111010000",
		"1001110111110000",
		"1001111000010000",
		"1001111000110001",
		"1001111001010001",
		"1001111001110010",
		"1001111010010010",
		"1001111010110011",
		"1001111011010011",
		"1001111011110100",
		"1001111100010101",
		"1001111100110110",
		"1001111101010111",
		"1001111101111000",
		"1001111110011001",
		"1001111110111010",
		"1001111111011011",
		"1001111111111100",
		"1010000000011110",
		"1010000000111111",
		"1010000001100000",
		"1010000010000010",
		"1010000010100011",
		"1010000011000101",
		"1010000011100110",
		"1010000100001000",
		"1010000100101010",
		"1010000101001100",
		"1010000101101101",
		"1010000110001111",
		"1010000110110001",
		"1010000111010011",
		"1010000111110101",
		"1010001000010111",
		"1010001000111010",
		"1010001001011100",
		"1010001001111110",
		"1010001010100001",
		"1010001011000011",
		"1010001011100101",
		"1010001100001000",
		"1010001100101010",
		"1010001101001101",
		"1010001101110000",
		"1010001110010011",
		"1010001110110101",
		"1010001111011000",
		"1010001111111011",
		"1010010000011110",
		"1010010001000001",
		"1010010001100100",
		"1010010010000111",
		"1010010010101010",
		"1010010011001110",
		"1010010011110001",
		"1010010100010100",
		"1010010100111000",
		"1010010101011011",
		"1010010101111111",
		"1010010110100010",
		"1010010111000110",
		"1010010111101010",
		"1010011000001101",
		"1010011000110001",
		"1010011001010101",
		"1010011001111001",
		"1010011010011101",
		"1010011011000001",
		"1010011011100101",
		"1010011100001001",
		"1010011100101101",
		"1010011101010001",
		"1010011101110110",
		"1010011110011010",
		"1010011110111110",
		"1010011111100011",
		"1010100000000111",
		"1010100000101100",
		"1010100001010000",
		"1010100001110101",
		"1010100010011010",
		"1010100010111110",
		"1010100011100011",
		"1010100100001000",
		"1010100100101101",
		"1010100101010010",
		"1010100101110111",
		"1010100110011100",
		"1010100111000001",
		"1010100111100110",
		"1010101000001100",
		"1010101000110001",
		"1010101001010110",
		"1010101001111011",
		"1010101010100001",
		"1010101011000110",
		"1010101011101100",
		"1010101100010001",
		"1010101100110111",
		"1010101101011101",
		"1010101110000011",
		"1010101110101000",
		"1010101111001110",
		"1010101111110100",
		"1010110000011010",
		"1010110001000000",
		"1010110001100110",
		"1010110010001100",
		"1010110010110010",
		"1010110011011000",
		"1010110011111111",
		"1010110100100101",
		"1010110101001011",
		"1010110101110010",
		"1010110110011000",
		"1010110110111111",
		"1010110111100101",
		"1010111000001100",
		"1010111000110010",
		"1010111001011001",
		"1010111010000000",
		"1010111010100111",
		"1010111011001101",
		"1010111011110100",
		"1010111100011011",
		"1010111101000010",
		"1010111101101001",
		"1010111110010000",
		"1010111110110111",
		"1010111111011111",
		"1011000000000110",
		"1011000000101101",
		"1011000001010100",
		"1011000001111100",
		"1011000010100011",
		"1011000011001011",
		"1011000011110010",
		"1011000100011010",
		"1011000101000001",
		"1011000101101001",
		"1011000110010001",
		"1011000110111000",
		"1011000111100000",
		"1011001000001000",
		"1011001000110000",
		"1011001001011000",
		"1011001010000000",
		"1011001010101000",
		"1011001011010000",
		"1011001011111000",
		"1011001100100000",
		"1011001101001000",
		"1011001101110001",
		"1011001110011001",
		"1011001111000001",
		"1011001111101010",
		"1011010000010010",
		"1011010000111011",
		"1011010001100011",
		"1011010010001100",
		"1011010010110100",
		"1011010011011101",
		"1011010100000110",
		"1011010100101110",
		"1011010101010111",
		"1011010110000000",
		"1011010110101001",
		"1011010111010010",
		"1011010111111011",
		"1011011000100100",
		"1011011001001101",
		"1011011001110110",
		"1011011010011111",
		"1011011011001000",
		"1011011011110010",
		"1011011100011011",
		"1011011101000100",
		"1011011101101110",
		"1011011110010111",
		"1011011111000001",
		"1011011111101010",
		"1011100000010100",
		"1011100000111101",
		"1011100001100111",
		"1011100010010001",
		"1011100010111010",
		"1011100011100100",
		"1011100100001110",
		"1011100100111000",
		"1011100101100010",
		"1011100110001100",
		"1011100110110110",
		"1011100111100000",
		"1011101000001010",
		"1011101000110100",
		"1011101001011110",
		"1011101010001000",
		"1011101010110010",
		"1011101011011101",
		"1011101100000111",
		"1011101100110001",
		"1011101101011100",
		"1011101110000110",
		"1011101110110001",
		"1011101111011011",
		"1011110000000110",
		"1011110000110000",
		"1011110001011011",
		"1011110010000110",
		"1011110010110000",
		"1011110011011011",
		"1011110100000110",
		"1011110100110001",
		"1011110101011100",
		"1011110110000111",
		"1011110110110010",
		"1011110111011101",
		"1011111000001000",
		"1011111000110011",
		"1011111001011110",
		"1011111010001001",
		"1011111010110100",
		"1011111011100000",
		"1011111100001011",
		"1011111100110110",
		"1011111101100010",
		"1011111110001101",
		"1011111110111001",
		"1011111111100100",
		"1100000000010000",
		"1100000000111011",
		"1100000001100111",
		"1100000010010010",
		"1100000010111110",
		"1100000011101010",
		"1100000100010101",
		"1100000101000001",
		"1100000101101101",
		"1100000110011001",
		"1100000111000101",
		"1100000111110001",
		"1100001000011101",
		"1100001001001001",
		"1100001001110101",
		"1100001010100001",
		"1100001011001101",
		"1100001011111001",
		"1100001100100101",
		"1100001101010010",
		"1100001101111110",
		"1100001110101010",
		"1100001111010111",
		"1100010000000011",
		"1100010000101111",
		"1100010001011100",
		"1100010010001000",
		"1100010010110101",
		"1100010011100001",
		"1100010100001110",
		"1100010100111011",
		"1100010101100111",
		"1100010110010100",
		"1100010111000001",
		"1100010111101110",
		"1100011000011010",
		"1100011001000111",
		"1100011001110100",
		"1100011010100001",
		"1100011011001110",
		"1100011011111011",
		"1100011100101000",
		"1100011101010101",
		"1100011110000010",
		"1100011110101111",
		"1100011111011100",
		"1100100000001010",
		"1100100000110111",
		"1100100001100100",
		"1100100010010001",
		"1100100010111111",
		"1100100011101100",
		"1100100100011001",
		"1100100101000111",
		"1100100101110100",
		"1100100110100010",
		"1100100111001111",
		"1100100111111101",
		"1100101000101010",
		"1100101001011000",
		"1100101010000110",
		"1100101010110011",
		"1100101011100001",
		"1100101100001111",
		"1100101100111101",
		"1100101101101010",
		"1100101110011000",
		"1100101111000110",
		"1100101111110100",
		"1100110000100010",
		"1100110001010000",
		"1100110001111110",
		"1100110010101100",
		"1100110011011010",
		"1100110100001000",
		"1100110100110110",
		"1100110101100100",
		"1100110110010011",
		"1100110111000001",
		"1100110111101111",
		"1100111000011101",
		"1100111001001100",
		"1100111001111010",
		"1100111010101000",
		"1100111011010111",
		"1100111100000101",
		"1100111100110100",
		"1100111101100010",
		"1100111110010001",
		"1100111110111111",
		"1100111111101110",
		"1101000000011100",
		"1101000001001011",
		"1101000001111010",
		"1101000010101000",
		"1101000011010111",
		"1101000100000110",
		"1101000100110100",
		"1101000101100011",
		"1101000110010010",
		"1101000111000001",
		"1101000111110000",
		"1101001000011111",
		"1101001001001110",
		"1101001001111101",
		"1101001010101100",
		"1101001011011011",
		"1101001100001010",
		"1101001100111001",
		"1101001101101000",
		"1101001110010111",
		"1101001111000110",
		"1101001111110101",
		"1101010000100101",
		"1101010001010100",
		"1101010010000011",
		"1101010010110010",
		"1101010011100010",
		"1101010100010001",
		"1101010101000000",
		"1101010101110000",
		"1101010110011111",
		"1101010111001111",
		"1101010111111110",
		"1101011000101110",
		"1101011001011101",
		"1101011010001101",
		"1101011010111100",
		"1101011011101100",
		"1101011100011011",
		"1101011101001011",
		"1101011101111011",
		"1101011110101010",
		"1101011111011010",
		"1101100000001010",
		"1101100000111010",
		"1101100001101001",
		"1101100010011001",
		"1101100011001001",
		"1101100011111001",
		"1101100100101001",
		"1101100101011001",
		"1101100110001001",
		"1101100110111001",
		"1101100111101001",
		"1101101000011001",
		"1101101001001001",
		"1101101001111001",
		"1101101010101001",
		"1101101011011001",
		"1101101100001001",
		"1101101100111001",
		"1101101101101001",
		"1101101110011001",
		"1101101111001010",
		"1101101111111010",
		"1101110000101010",
		"1101110001011010",
		"1101110010001011",
		"1101110010111011",
		"1101110011101011",
		"1101110100011100",
		"1101110101001100",
		"1101110101111100",
		"1101110110101101",
		"1101110111011101",
		"1101111000001110",
		"1101111000111110",
		"1101111001101111",
		"1101111010011111",
		"1101111011010000",
		"1101111100000000",
		"1101111100110001",
		"1101111101100001",
		"1101111110010010",
		"1101111111000011",
		"1101111111110011",
		"1110000000100100",
		"1110000001010101",
		"1110000010000101",
		"1110000010110110",
		"1110000011100111",
		"1110000100011000",
		"1110000101001000",
		"1110000101111001",
		"1110000110101010",
		"1110000111011011",
		"1110001000001100",
		"1110001000111101",
		"1110001001101101",
		"1110001010011110",
		"1110001011001111",
		"1110001100000000",
		"1110001100110001",
		"1110001101100010",
		"1110001110010011",
		"1110001111000100",
		"1110001111110101",
		"1110010000100110",
		"1110010001010111",
		"1110010010001000",
		"1110010010111010",
		"1110010011101011",
		"1110010100011100",
		"1110010101001101",
		"1110010101111110",
		"1110010110101111",
		"1110010111100000",
		"1110011000010010",
		"1110011001000011",
		"1110011001110100",
		"1110011010100101",
		"1110011011010111",
		"1110011100001000",
		"1110011100111001",
		"1110011101101011",
		"1110011110011100",
		"1110011111001101",
		"1110011111111111",
		"1110100000110000",
		"1110100001100001",
		"1110100010010011",
		"1110100011000100",
		"1110100011110110",
		"1110100100100111",
		"1110100101011001",
		"1110100110001010",
		"1110100110111100",
		"1110100111101101",
		"1110101000011111",
		"1110101001010000",
		"1110101010000010",
		"1110101010110011",
		"1110101011100101",
		"1110101100010110",
		"1110101101001000",
		"1110101101111010",
		"1110101110101011",
		"1110101111011101",
		"1110110000001110",
		"1110110001000000",
		"1110110001110010",
		"1110110010100011",
		"1110110011010101",
		"1110110100000111",
		"1110110100111001",
		"1110110101101010",
		"1110110110011100",
		"1110110111001110",
		"1110111000000000",
		"1110111000110001",
		"1110111001100011",
		"1110111010010101",
		"1110111011000111",
		"1110111011111001",
		"1110111100101010",
		"1110111101011100",
		"1110111110001110",
		"1110111111000000",
		"1110111111110010",
		"1111000000100100",
		"1111000001010101",
		"1111000010000111",
		"1111000010111001",
		"1111000011101011",
		"1111000100011101",
		"1111000101001111",
		"1111000110000001",
		"1111000110110011",
		"1111000111100101",
		"1111001000010111",
		"1111001001001001",
		"1111001001111011",
		"1111001010101101",
		"1111001011011111",
		"1111001100010001",
		"1111001101000011",
		"1111001101110101",
		"1111001110100111",
		"1111001111011001",
		"1111010000001011",
		"1111010000111101",
		"1111010001101111",
		"1111010010100001",
		"1111010011010011",
		"1111010100000101",
		"1111010100110111",
		"1111010101101001",
		"1111010110011011",
		"1111010111001110",
		"1111011000000000",
		"1111011000110010",
		"1111011001100100",
		"1111011010010110",
		"1111011011001000",
		"1111011011111010",
		"1111011100101100",
		"1111011101011111",
		"1111011110010001",
		"1111011111000011",
		"1111011111110101",
		"1111100000100111",
		"1111100001011001",
		"1111100010001100",
		"1111100010111110",
		"1111100011110000",
		"1111100100100010",
		"1111100101010100",
		"1111100110000110",
		"1111100110111001",
		"1111100111101011",
		"1111101000011101",
		"1111101001001111",
		"1111101010000010",
		"1111101010110100",
		"1111101011100110",
		"1111101100011000",
		"1111101101001010",
		"1111101101111101",
		"1111101110101111",
		"1111101111100001",
		"1111110000010011",
		"1111110001000110",
		"1111110001111000",
		"1111110010101010",
		"1111110011011100",
		"1111110100001111",
		"1111110101000001",
		"1111110101110011",
		"1111110110100101",
		"1111110111011000",
		"1111111000001010",
		"1111111000111100",
		"1111111001101110",
		"1111111010100001",
		"1111111011010011",
		"1111111100000101",
		"1111111100110111",
		"1111111101101010",
		"1111111110011100",
		"1111111111001110",
		"0000000000000000",
		"0000000000110010",
		"0000000001100100",
		"0000000010010110",
		"0000000011001001",
		"0000000011111011",
		"0000000100101101",
		"0000000101011111",
		"0000000110010010",
		"0000000111000100",
		"0000000111110110",
		"0000001000101000",
		"0000001001011011",
		"0000001010001101",
		"0000001010111111",
		"0000001011110001",
		"0000001100100100",
		"0000001101010110",
		"0000001110001000",
		"0000001110111010",
		"0000001111101101",
		"0000010000011111",
		"0000010001010001",
		"0000010010000011",
		"0000010010110110",
		"0000010011101000",
		"0000010100011010",
		"0000010101001100",
		"0000010101111110",
		"0000010110110001",
		"0000010111100011",
		"0000011000010101",
		"0000011001000111",
		"0000011001111010",
		"0000011010101100",
		"0000011011011110",
		"0000011100010000",
		"0000011101000010",
		"0000011101110100",
		"0000011110100111",
		"0000011111011001",
		"0000100000001011",
		"0000100000111101",
		"0000100001101111",
		"0000100010100001",
		"0000100011010100",
		"0000100100000110",
		"0000100100111000",
		"0000100101101010",
		"0000100110011100",
		"0000100111001110",
		"0000101000000000",
		"0000101000110010",
		"0000101001100101",
		"0000101010010111",
		"0000101011001001",
		"0000101011111011",
		"0000101100101101",
		"0000101101011111",
		"0000101110010001",
		"0000101111000011",
		"0000101111110101",
		"0000110000100111",
		"0000110001011001",
		"0000110010001011",
		"0000110010111101",
		"0000110011101111",
		"0000110100100001",
		"0000110101010011",
		"0000110110000101",
		"0000110110110111",
		"0000110111101001",
		"0000111000011011",
		"0000111001001101",
		"0000111001111111",
		"0000111010110001",
		"0000111011100011",
		"0000111100010101",
		"0000111101000111",
		"0000111101111001",
		"0000111110101011",
		"0000111111011100",
		"0001000000001110",
		"0001000001000000",
		"0001000001110010",
		"0001000010100100",
		"0001000011010110",
		"0001000100000111",
		"0001000100111001",
		"0001000101101011",
		"0001000110011101",
		"0001000111001111",
		"0001001000000000",
		"0001001000110010",
		"0001001001100100",
		"0001001010010110",
		"0001001011000111",
		"0001001011111001",
		"0001001100101011",
		"0001001101011101",
		"0001001110001110",
		"0001001111000000",
		"0001001111110010",
		"0001010000100011",
		"0001010001010101",
		"0001010010000110",
		"0001010010111000",
		"0001010011101010",
		"0001010100011011",
		"0001010101001101",
		"0001010101111110",
		"0001010110110000",
		"0001010111100001",
		"0001011000010011",
		"0001011001000100",
		"0001011001110110",
		"0001011010100111",
		"0001011011011001",
		"0001011100001010",
		"0001011100111100",
		"0001011101101101",
		"0001011110011111",
		"0001011111010000",
		"0001100000000001",
		"0001100000110011",
		"0001100001100100",
		"0001100010010101",
		"0001100011000111",
		"0001100011111000",
		"0001100100101001",
		"0001100101011011",
		"0001100110001100",
		"0001100110111101",
		"0001100111101110",
		"0001101000100000",
		"0001101001010001",
		"0001101010000010",
		"0001101010110011",
		"0001101011100100",
		"0001101100010101",
		"0001101101000110",
		"0001101101111000",
		"0001101110101001",
		"0001101111011010",
		"0001110000001011",
		"0001110000111100",
		"0001110001101101",
		"0001110010011110",
		"0001110011001111",
		"0001110100000000",
		"0001110100110001",
		"0001110101100010",
		"0001110110010011",
		"0001110111000011",
		"0001110111110100",
		"0001111000100101",
		"0001111001010110",
		"0001111010000111",
		"0001111010111000",
		"0001111011101000",
		"0001111100011001",
		"0001111101001010",
		"0001111101111011",
		"0001111110101011",
		"0001111111011100",
		"0010000000001101",
		"0010000000111101",
		"0010000001101110",
		"0010000010011111",
		"0010000011001111",
		"0010000100000000",
		"0010000100110000",
		"0010000101100001",
		"0010000110010001",
		"0010000111000010",
		"0010000111110010",
		"0010001000100011",
		"0010001001010011",
		"0010001010000100",
		"0010001010110100",
		"0010001011100100",
		"0010001100010101",
		"0010001101000101",
		"0010001101110101",
		"0010001110100110",
		"0010001111010110",
		"0010010000000110",
		"0010010000110110",
		"0010010001100111",
		"0010010010010111",
		"0010010011000111",
		"0010010011110111",
		"0010010100100111",
		"0010010101010111",
		"0010010110000111",
		"0010010110110111",
		"0010010111100111",
		"0010011000010111",
		"0010011001000111",
		"0010011001110111",
		"0010011010100111",
		"0010011011010111",
		"0010011100000111",
		"0010011100110111",
		"0010011101100111",
		"0010011110010111",
		"0010011111000110",
		"0010011111110110",
		"0010100000100110",
		"0010100001010110",
		"0010100010000101",
		"0010100010110101",
		"0010100011100101",
		"0010100100010100",
		"0010100101000100",
		"0010100101110011",
		"0010100110100011",
		"0010100111010010",
		"0010101000000010",
		"0010101000110001",
		"0010101001100001",
		"0010101010010000",
		"0010101011000000",
		"0010101011101111",
		"0010101100011110",
		"0010101101001110",
		"0010101101111101",
		"0010101110101100",
		"0010101111011011",
		"0010110000001011",
		"0010110000111010",
		"0010110001101001",
		"0010110010011000",
		"0010110011000111",
		"0010110011110110",
		"0010110100100101",
		"0010110101010100",
		"0010110110000011",
		"0010110110110010",
		"0010110111100001",
		"0010111000010000",
		"0010111000111111",
		"0010111001101110",
		"0010111010011101",
		"0010111011001100",
		"0010111011111010",
		"0010111100101001",
		"0010111101011000",
		"0010111110000110",
		"0010111110110101",
		"0010111111100100",
		"0011000000010010",
		"0011000001000001",
		"0011000001101111",
		"0011000010011110",
		"0011000011001100",
		"0011000011111011",
		"0011000100101001",
		"0011000101011000",
		"0011000110000110",
		"0011000110110100",
		"0011000111100011",
		"0011001000010001",
		"0011001000111111",
		"0011001001101101",
		"0011001010011100",
		"0011001011001010",
		"0011001011111000",
		"0011001100100110",
		"0011001101010100",
		"0011001110000010",
		"0011001110110000",
		"0011001111011110",
		"0011010000001100",
		"0011010000111010",
		"0011010001101000",
		"0011010010010110",
		"0011010011000011",
		"0011010011110001",
		"0011010100011111",
		"0011010101001101",
		"0011010101111010",
		"0011010110101000",
		"0011010111010110",
		"0011011000000011",
		"0011011000110001",
		"0011011001011110",
		"0011011010001100",
		"0011011010111001",
		"0011011011100111",
		"0011011100010100",
		"0011011101000001",
		"0011011101101111",
		"0011011110011100",
		"0011011111001001",
		"0011011111110110",
		"0011100000100100",
		"0011100001010001",
		"0011100001111110",
		"0011100010101011",
		"0011100011011000",
		"0011100100000101",
		"0011100100110010",
		"0011100101011111",
		"0011100110001100",
		"0011100110111001",
		"0011100111100110",
		"0011101000010010",
		"0011101000111111",
		"0011101001101100",
		"0011101010011001",
		"0011101011000101",
		"0011101011110010",
		"0011101100011111",
		"0011101101001011",
		"0011101101111000",
		"0011101110100100",
		"0011101111010001",
		"0011101111111101",
		"0011110000101001",
		"0011110001010110",
		"0011110010000010",
		"0011110010101110",
		"0011110011011011",
		"0011110100000111",
		"0011110100110011",
		"0011110101011111",
		"0011110110001011",
		"0011110110110111",
		"0011110111100011",
		"0011111000001111",
		"0011111000111011",
		"0011111001100111",
		"0011111010010011",
		"0011111010111111",
		"0011111011101011",
		"0011111100010110",
		"0011111101000010",
		"0011111101101110",
		"0011111110011001",
		"0011111111000101",
		"0011111111110000",
		"0100000000011100",
		"0100000001000111",
		"0100000001110011",
		"0100000010011110",
		"0100000011001010",
		"0100000011110101",
		"0100000100100000",
		"0100000101001100",
		"0100000101110111",
		"0100000110100010",
		"0100000111001101",
		"0100000111111000",
		"0100001000100011",
		"0100001001001110",
		"0100001001111001",
		"0100001010100100",
		"0100001011001111",
		"0100001011111010",
		"0100001100100101",
		"0100001101010000",
		"0100001101111010",
		"0100001110100101",
		"0100001111010000",
		"0100001111111010",
		"0100010000100101",
		"0100010001001111",
		"0100010001111010",
		"0100010010100100",
		"0100010011001111",
		"0100010011111001",
		"0100010100100011",
		"0100010101001110",
		"0100010101111000",
		"0100010110100010",
		"0100010111001100",
		"0100010111110110",
		"0100011000100000",
		"0100011001001010",
		"0100011001110100",
		"0100011010011110",
		"0100011011001000",
		"0100011011110010",
		"0100011100011100",
		"0100011101000110",
		"0100011101101111",
		"0100011110011001",
		"0100011111000011",
		"0100011111101100",
		"0100100000010110",
		"0100100000111111",
		"0100100001101001",
		"0100100010010010",
		"0100100010111100",
		"0100100011100101",
		"0100100100001110",
		"0100100100111000",
		"0100100101100001",
		"0100100110001010",
		"0100100110110011",
		"0100100111011100",
		"0100101000000101",
		"0100101000101110",
		"0100101001010111",
		"0100101010000000",
		"0100101010101001",
		"0100101011010010",
		"0100101011111010",
		"0100101100100011",
		"0100101101001100",
		"0100101101110100",
		"0100101110011101",
		"0100101111000101",
		"0100101111101110",
		"0100110000010110",
		"0100110000111111",
		"0100110001100111",
		"0100110010001111",
		"0100110010111000",
		"0100110011100000",
		"0100110100001000",
		"0100110100110000",
		"0100110101011000",
		"0100110110000000",
		"0100110110101000",
		"0100110111010000",
		"0100110111111000",
		"0100111000100000",
		"0100111001001000",
		"0100111001101111",
		"0100111010010111",
		"0100111010111111",
		"0100111011100110",
		"0100111100001110",
		"0100111100110101",
		"0100111101011101",
		"0100111110000100",
		"0100111110101100",
		"0100111111010011",
		"0100111111111010",
		"0101000000100001",
		"0101000001001001",
		"0101000001110000",
		"0101000010010111",
		"0101000010111110",
		"0101000011100101",
		"0101000100001100",
		"0101000100110011",
		"0101000101011001",
		"0101000110000000",
		"0101000110100111",
		"0101000111001110",
		"0101000111110100",
		"0101001000011011",
		"0101001001000001",
		"0101001001101000",
		"0101001010001110",
		"0101001010110101",
		"0101001011011011",
		"0101001100000001",
		"0101001100101000",
		"0101001101001110",
		"0101001101110100",
		"0101001110011010",
		"0101001111000000",
		"0101001111100110",
		"0101010000001100",
		"0101010000110010",
		"0101010001011000",
		"0101010001111101",
		"0101010010100011",
		"0101010011001001",
		"0101010011101111",
		"0101010100010100",
		"0101010100111010",
		"0101010101011111",
		"0101010110000101",
		"0101010110101010",
		"0101010111001111",
		"0101010111110100",
		"0101011000011010",
		"0101011000111111",
		"0101011001100100",
		"0101011010001001",
		"0101011010101110",
		"0101011011010011",
		"0101011011111000",
		"0101011100011101",
		"0101011101000010",
		"0101011101100110",
		"0101011110001011",
		"0101011110110000",
		"0101011111010100",
		"0101011111111001",
		"0101100000011101",
		"0101100001000010",
		"0101100001100110",
		"0101100010001010",
		"0101100010101111",
		"0101100011010011",
		"0101100011110111",
		"0101100100011011",
		"0101100100111111",
		"0101100101100011",
		"0101100110000111",
		"0101100110101011",
		"0101100111001111",
		"0101100111110011",
		"0101101000010110",
		"0101101000111010",
		"0101101001011110",
		"0101101010000001",
		"0101101010100101",
		"0101101011001000",
		"0101101011101100",
		"0101101100001111",
		"0101101100110010",
		"0101101101010110",
		"0101101101111001",
		"0101101110011100",
		"0101101110111111",
		"0101101111100010",
		"0101110000000101",
		"0101110000101000",
		"0101110001001011",
		"0101110001101101",
		"0101110010010000",
		"0101110010110011",
		"0101110011010110",
		"0101110011111000",
		"0101110100011011",
		"0101110100111101",
		"0101110101011111",
		"0101110110000010",
		"0101110110100100",
		"0101110111000110",
		"0101110111101001",
		"0101111000001011",
		"0101111000101101",
		"0101111001001111",
		"0101111001110001",
		"0101111010010011",
		"0101111010110100",
		"0101111011010110",
		"0101111011111000",
		"0101111100011010",
		"0101111100111011",
		"0101111101011101",
		"0101111101111110",
		"0101111110100000",
		"0101111111000001",
		"0101111111100010",
		"0110000000000100",
		"0110000000100101",
		"0110000001000110",
		"0110000001100111",
		"0110000010001000",
		"0110000010101001",
		"0110000011001010",
		"0110000011101011",
		"0110000100001100",
		"0110000100101101",
		"0110000101001101",
		"0110000101101110",
		"0110000110001110",
		"0110000110101111",
		"0110000111001111",
		"0110000111110000",
		"0110001000010000",
		"0110001000110000",
		"0110001001010001",
		"0110001001110001",
		"0110001010010001",
		"0110001010110001",
		"0110001011010001",
		"0110001011110001",
		"0110001100010001",
		"0110001100110000",
		"0110001101010000",
		"0110001101110000",
		"0110001110001111",
		"0110001110101111",
		"0110001111001110",
		"0110001111101110",
		"0110010000001101",
		"0110010000101101",
		"0110010001001100",
		"0110010001101011",
		"0110010010001010",
		"0110010010101001",
		"0110010011001000",
		"0110010011100111",
		"0110010100000110",
		"0110010100100101",
		"0110010101000100",
		"0110010101100010",
		"0110010110000001",
		"0110010110100000",
		"0110010110111110",
		"0110010111011101",
		"0110010111111011",
		"0110011000011001",
		"0110011000111000",
		"0110011001010110",
		"0110011001110100",
		"0110011010010010",
		"0110011010110000",
		"0110011011001110",
		"0110011011101100",
		"0110011100001010",
		"0110011100101000",
		"0110011101000101",
		"0110011101100011",
		"0110011110000001",
		"0110011110011110",
		"0110011110111100",
		"0110011111011001",
		"0110011111110111",
		"0110100000010100",
		"0110100000110001",
		"0110100001001110",
		"0110100001101011",
		"0110100010001000",
		"0110100010100101",
		"0110100011000010",
		"0110100011011111",
		"0110100011111100",
		"0110100100011001",
		"0110100100110101",
		"0110100101010010",
		"0110100101101110",
		"0110100110001011",
		"0110100110100111",
		"0110100111000100",
		"0110100111100000",
		"0110100111111100",
		"0110101000011000",
		"0110101000110100",
		"0110101001010000",
		"0110101001101100",
		"0110101010001000",
		"0110101010100100",
		"0110101011000000",
		"0110101011011011",
		"0110101011110111",
		"0110101100010011",
		"0110101100101110",
		"0110101101001010",
		"0110101101100101",
		"0110101110000000",
		"0110101110011100",
		"0110101110110111",
		"0110101111010010",
		"0110101111101101",
		"0110110000001000",
		"0110110000100011",
		"0110110000111110",
		"0110110001011000",
		"0110110001110011",
		"0110110010001110",
		"0110110010101000",
		"0110110011000011",
		"0110110011011101",
		"0110110011111000",
		"0110110100010010",
		"0110110100101100",
		"0110110101000111",
		"0110110101100001",
		"0110110101111011",
		"0110110110010101",
		"0110110110101111",
		"0110110111001001",
		"0110110111100011",
		"0110110111111100",
		"0110111000010110",
		"0110111000110000",
		"0110111001001001",
		"0110111001100011",
		"0110111001111100",
		"0110111010010101",
		"0110111010101111",
		"0110111011001000",
		"0110111011100001",
		"0110111011111010",
		"0110111100010011",
		"0110111100101100",
		"0110111101000101",
		"0110111101011110",
		"0110111101110110",
		"0110111110001111",
		"0110111110101000",
		"0110111111000000",
		"0110111111011001",
		"0110111111110001",
		"0111000000001001",
		"0111000000100010",
		"0111000000111010",
		"0111000001010010",
		"0111000001101010",
		"0111000010000010",
		"0111000010011010",
		"0111000010110010",
		"0111000011001010",
		"0111000011100001",
		"0111000011111001",
		"0111000100010001",
		"0111000100101000",
		"0111000101000000",
		"0111000101010111",
		"0111000101101110",
		"0111000110000110",
		"0111000110011101",
		"0111000110110100",
		"0111000111001011",
		"0111000111100010",
		"0111000111111001",
		"0111001000010000",
		"0111001000100110",
		"0111001000111101",
		"0111001001010100",
		"0111001001101010",
		"0111001010000001",
		"0111001010010111",
		"0111001010101110",
		"0111001011000100",
		"0111001011011010",
		"0111001011110000",
		"0111001100000110",
		"0111001100011100",
		"0111001100110010",
		"0111001101001000",
		"0111001101011110",
		"0111001101110100",
		"0111001110001001",
		"0111001110011111",
		"0111001110110101",
		"0111001111001010",
		"0111001111011111",
		"0111001111110101",
		"0111010000001010",
		"0111010000011111",
		"0111010000110100",
		"0111010001001001",
		"0111010001011110",
		"0111010001110011",
		"0111010010001000",
		"0111010010011101",
		"0111010010110001",
		"0111010011000110",
		"0111010011011011",
		"0111010011101111",
		"0111010100000011",
		"0111010100011000",
		"0111010100101100",
		"0111010101000000",
		"0111010101010100",
		"0111010101101000",
		"0111010101111100",
		"0111010110010000",
		"0111010110100100",
		"0111010110111000",
		"0111010111001100",
		"0111010111011111",
		"0111010111110011",
		"0111011000000110",
		"0111011000011010",
		"0111011000101101",
		"0111011001000000",
		"0111011001010011",
		"0111011001100111",
		"0111011001111010",
		"0111011010001101",
		"0111011010100000",
		"0111011010110010",
		"0111011011000101",
		"0111011011011000",
		"0111011011101010",
		"0111011011111101",
		"0111011100010000",
		"0111011100100010",
		"0111011100110100",
		"0111011101000111",
		"0111011101011001",
		"0111011101101011",
		"0111011101111101",
		"0111011110001111",
		"0111011110100001",
		"0111011110110011",
		"0111011111000100",
		"0111011111010110",
		"0111011111101000",
		"0111011111111001",
		"0111100000001011",
		"0111100000011100",
		"0111100000101110",
		"0111100000111111",
		"0111100001010000",
		"0111100001100001",
		"0111100001110010",
		"0111100010000011",
		"0111100010010100",
		"0111100010100101",
		"0111100010110110",
		"0111100011000110",
		"0111100011010111",
		"0111100011100111",
		"0111100011111000",
		"0111100100001000",
		"0111100100011001",
		"0111100100101001",
		"0111100100111001",
		"0111100101001001",
		"0111100101011001",
		"0111100101101001",
		"0111100101111001",
		"0111100110001001",
		"0111100110011000",
		"0111100110101000",
		"0111100110111000",
		"0111100111000111",
		"0111100111010111",
		"0111100111100110",
		"0111100111110101",
		"0111101000000100",
		"0111101000010100",
		"0111101000100011",
		"0111101000110010",
		"0111101001000001",
		"0111101001001111",
		"0111101001011110",
		"0111101001101101",
		"0111101001111100",
		"0111101010001010",
		"0111101010011001",
		"0111101010100111",
		"0111101010110101",
		"0111101011000100",
		"0111101011010010",
		"0111101011100000",
		"0111101011101110",
		"0111101011111100",
		"0111101100001010",
		"0111101100011000",
		"0111101100100101",
		"0111101100110011",
		"0111101101000001",
		"0111101101001110",
		"0111101101011100",
		"0111101101101001",
		"0111101101110110",
		"0111101110000011",
		"0111101110010001",
		"0111101110011110",
		"0111101110101011",
		"0111101110111000",
		"0111101111000100",
		"0111101111010001",
		"0111101111011110",
		"0111101111101011",
		"0111101111110111",
		"0111110000000100",
		"0111110000010000",
		"0111110000011100",
		"0111110000101001",
		"0111110000110101",
		"0111110001000001",
		"0111110001001101",
		"0111110001011001",
		"0111110001100101",
		"0111110001110000",
		"0111110001111100",
		"0111110010001000",
		"0111110010010011",
		"0111110010011111",
		"0111110010101010",
		"0111110010110110",
		"0111110011000001",
		"0111110011001100",
		"0111110011010111",
		"0111110011100010",
		"0111110011101101",
		"0111110011111000",
		"0111110100000011",
		"0111110100001110",
		"0111110100011000",
		"0111110100100011",
		"0111110100101110",
		"0111110100111000",
		"0111110101000010",
		"0111110101001101",
		"0111110101010111",
		"0111110101100001",
		"0111110101101011",
		"0111110101110101",
		"0111110101111111",
		"0111110110001001",
		"0111110110010011",
		"0111110110011100",
		"0111110110100110",
		"0111110110110000",
		"0111110110111001",
		"0111110111000010",
		"0111110111001100",
		"0111110111010101",
		"0111110111011110",
		"0111110111100111",
		"0111110111110000",
		"0111110111111001",
		"0111111000000010",
		"0111111000001011",
		"0111111000010011",
		"0111111000011100",
		"0111111000100101",
		"0111111000101101",
		"0111111000110110",
		"0111111000111110",
		"0111111001000110",
		"0111111001001110",
		"0111111001010110",
		"0111111001011110",
		"0111111001100110",
		"0111111001101110",
		"0111111001110110",
		"0111111001111110",
		"0111111010000101",
		"0111111010001101",
		"0111111010010100",
		"0111111010011100",
		"0111111010100011",
		"0111111010101010",
		"0111111010110010",
		"0111111010111001",
		"0111111011000000",
		"0111111011000111",
		"0111111011001110",
		"0111111011010100",
		"0111111011011011",
		"0111111011100010",
		"0111111011101000",
		"0111111011101111",
		"0111111011110101",
		"0111111011111100",
		"0111111100000010",
		"0111111100001000",
		"0111111100001110",
		"0111111100010100",
		"0111111100011010",
		"0111111100100000",
		"0111111100100110",
		"0111111100101100",
		"0111111100110001",
		"0111111100110111",
		"0111111100111100",
		"0111111101000010",
		"0111111101000111",
		"0111111101001100",
		"0111111101010010",
		"0111111101010111",
		"0111111101011100",
		"0111111101100001",
		"0111111101100110",
		"0111111101101010",
		"0111111101101111",
		"0111111101110100",
		"0111111101111000",
		"0111111101111101",
		"0111111110000001",
		"0111111110000110",
		"0111111110001010",
		"0111111110001110",
		"0111111110010010",
		"0111111110010110",
		"0111111110011010",
		"0111111110011110",
		"0111111110100010",
		"0111111110100110",
		"0111111110101001",
		"0111111110101101",
		"0111111110110000",
		"0111111110110100",
		"0111111110110111",
		"0111111110111011",
		"0111111110111110",
		"0111111111000001",
		"0111111111000100",
		"0111111111000111",
		"0111111111001010",
		"0111111111001101",
		"0111111111001111",
		"0111111111010010",
		"0111111111010101",
		"0111111111010111",
		"0111111111011001",
		"0111111111011100",
		"0111111111011110",
		"0111111111100000",
		"0111111111100010",
		"0111111111100100",
		"0111111111100110",
		"0111111111101000",
		"0111111111101010",
		"0111111111101100",
		"0111111111101110",
		"0111111111101111",
		"0111111111110001",
		"0111111111110010",
		"0111111111110011",
		"0111111111110101",
		"0111111111110110",
		"0111111111110111",
		"0111111111111000",
		"0111111111111001",
		"0111111111111010",
		"0111111111111011",
		"0111111111111011",
		"0111111111111100",
		"0111111111111101",
		"0111111111111101",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110",
		"0111111111111110");
begin

	process(clk)
	begin
		if rising_edge(clk) then
			data_a<=my_rom(to_integer(unsigned(addr_a)));
		end if;
	end process;
	process(clk)
	begin
		if rising_edge(clk) then
			data_b<=my_rom(to_integer(unsigned(addr_b)));
		end if;
	end process;
end architecture behavioral;
